module andGate(a,b,and_out);
input a,b;
output and_out;

assign and_out = a & b;

endmodule