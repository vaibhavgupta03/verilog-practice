module halfAdder(
    input a,
    input b,
    output sum,
    output carry
);
    assign sum = a ^ b;      // Sum is the XOR of a and b
    assign carry = a & b;    // Carry is the AND of a and b
endmodule